
module InstructionMemory(Address, Instruction);
	input [31:0] Address;
	output reg [31:0] Instruction;
	
	always @(*)
		case (Address[9:2])//pay attention to j,jal, in MARS the PC begin at 0x00400000 but in our CPU it's 0x0
		
			8'd0: Instruction<=32'h08100003;
			8'd1: Instruction<=32'h08100028;
			8'd2: Instruction<=32'h0810008b;
			8'd3: Instruction<=32'h3c044000;
			8'd4: Instruction<=32'h20050000;
			8'd5: Instruction<=32'h20060000;
			8'd6: Instruction<=32'h20070000;
			8'd7: Instruction<=32'h200c0001;
			8'd8: Instruction<=32'h200d0002;
			8'd9: Instruction<=32'h200e0003;
			8'd10: Instruction<=32'h200ffff9;
			8'd11: Instruction<=32'h2018ffff;
			8'd12: Instruction<=32'h8c910014;
			8'd13: Instruction<=32'h00000000;
			8'd14: Instruction<=32'h00000000;
			8'd15: Instruction<=32'h00000000;
			8'd16: Instruction<=32'h00000000;
			8'd17: Instruction<=32'h00000000;
			8'd18: Instruction<=32'h00000000;
			8'd19: Instruction<=32'h00000000;
			8'd20: Instruction<=32'h00000000;
			8'd21: Instruction<=32'h00000000;
			8'd22: Instruction<=32'h00000000;
			8'd23: Instruction<=32'h00000000;
			8'd24: Instruction<=32'h00000000;
			8'd25: Instruction<=32'h00000000;
			8'd26: Instruction<=32'h00000000;
			8'd27: Instruction<=32'h00000000;
			8'd28: Instruction<=32'h00000000;
			8'd29: Instruction<=32'h00000000;
			8'd30: Instruction<=32'h00000000;
			8'd31: Instruction<=32'h00000000;
			8'd32: Instruction<=32'h00000000;
			8'd33: Instruction<=32'h8c920014;
			8'd34: Instruction<=32'h02513022;
			8'd35: Instruction<=32'h2010fffb;
			8'd36: Instruction<=32'hac900000;
			8'd37: Instruction<=32'hac980004;
			8'd38: Instruction<=32'hac8e0008;
			8'd39: Instruction<=32'h0810008c;
			8'd40: Instruction<=32'h8c880008;
			8'd41: Instruction<=32'h010f4024;
			8'd42: Instruction<=32'hac880008;
			8'd43: Instruction<=32'h10a0000b;
			8'd44: Instruction<=32'h10ac000e;
			8'd45: Instruction<=32'h10ad0012;
			8'd46: Instruction<=32'h10ae0016;
			8'd47: Instruction<=32'hac870010;
			8'd48: Instruction<=32'h14ae0001;
			8'd49: Instruction<=32'h2005ffff;
			8'd50: Instruction<=32'h20a50001;
			8'd51: Instruction<=32'h8c880008;
			8'd52: Instruction<=32'h35080002;
			8'd53: Instruction<=32'hac880008;
			8'd54: Instruction<=32'h03400008;
			8'd55: Instruction<=32'h30d5000f;
			8'd56: Instruction<=32'h0c10004a;
			8'd57: Instruction<=32'h20e70100;
			8'd58: Instruction<=32'h0810002f;
			8'd59: Instruction<=32'h30d500f0;
			8'd60: Instruction<=32'h0015a902;
			8'd61: Instruction<=32'h0c10004a;
			8'd62: Instruction<=32'h20e70200;
			8'd63: Instruction<=32'h0810002f;
			8'd64: Instruction<=32'h30d50f00;
			8'd65: Instruction<=32'h0015aa02;
			8'd66: Instruction<=32'h0c10004a;
			8'd67: Instruction<=32'h20e70400;
			8'd68: Instruction<=32'h0810002f;
			8'd69: Instruction<=32'h30d5f000;
			8'd70: Instruction<=32'h0015ac02;
			8'd71: Instruction<=32'h0c10004a;
			8'd72: Instruction<=32'h20e70800;
			8'd73: Instruction<=32'h0810002f;
			8'd74: Instruction<=32'h20070000;
			8'd75: Instruction<=32'h22a80000;
			8'd76: Instruction<=32'h1100001e;
			8'd77: Instruction<=32'h22a8ffff;
			8'd78: Instruction<=32'h1100001e;
			8'd79: Instruction<=32'h22a8fffe;
			8'd80: Instruction<=32'h1100001e;
			8'd81: Instruction<=32'h22a8fffd;
			8'd82: Instruction<=32'h1100001e;
			8'd83: Instruction<=32'h22a8fffc;
			8'd84: Instruction<=32'h1100001e;
			8'd85: Instruction<=32'h22a8fffb;
			8'd86: Instruction<=32'h1100001e;
			8'd87: Instruction<=32'h22a8fffa;
			8'd88: Instruction<=32'h1100001e;
			8'd89: Instruction<=32'h22a8fff9;
			8'd90: Instruction<=32'h1100001e;
			8'd91: Instruction<=32'h22a8fff8;
			8'd92: Instruction<=32'h1100001e;
			8'd93: Instruction<=32'h22a8fff7;
			8'd94: Instruction<=32'h1100001e;
			8'd95: Instruction<=32'h22a8fff6;
			8'd96: Instruction<=32'h1100001e;
			8'd97: Instruction<=32'h22a8fff5;
			8'd98: Instruction<=32'h1100001e;
			8'd99: Instruction<=32'h22a8fff4;
			8'd100: Instruction<=32'h1100001e;
			8'd101: Instruction<=32'h22a8fff3;
			8'd102: Instruction<=32'h1100001e;
			8'd103: Instruction<=32'h22a8fff2;
			8'd104: Instruction<=32'h1100001e;
			8'd105: Instruction<=32'h22a8fff1;
			8'd106: Instruction<=32'h1100001e;
			8'd107: Instruction<=32'h2007003f;
			8'd108: Instruction<=32'h03e00008;
			8'd109: Instruction<=32'h20070006;
			8'd110: Instruction<=32'h03e00008;
			8'd111: Instruction<=32'h2007005b;
			8'd112: Instruction<=32'h03e00008;
			8'd113: Instruction<=32'h2007004f;
			8'd114: Instruction<=32'h03e00008;
			8'd115: Instruction<=32'h20070066;
			8'd116: Instruction<=32'h03e00008;
			8'd117: Instruction<=32'h2007006d;
			8'd118: Instruction<=32'h03e00008;
			8'd119: Instruction<=32'h2007007d;
			8'd120: Instruction<=32'h03e00008;
			8'd121: Instruction<=32'h20070007;
			8'd122: Instruction<=32'h03e00008;
			8'd123: Instruction<=32'h2007007f;
			8'd124: Instruction<=32'h03e00008;
			8'd125: Instruction<=32'h2007006f;
			8'd126: Instruction<=32'h03e00008;
			8'd127: Instruction<=32'h20070077;
			8'd128: Instruction<=32'h03e00008;
			8'd129: Instruction<=32'h2007007c;
			8'd130: Instruction<=32'h03e00008;
			8'd131: Instruction<=32'h20070039;
			8'd132: Instruction<=32'h03e00008;
			8'd133: Instruction<=32'h2007005e;
			8'd134: Instruction<=32'h03e00008;
			8'd135: Instruction<=32'h20070079;
			8'd136: Instruction<=32'h03e00008;
			8'd137: Instruction<=32'h20070071;
			8'd138: Instruction<=32'h03e00008;
			8'd139: Instruction<=32'h03400008;
			8'd140: Instruction<=32'h00000000;
			
			default: Instruction <= 32'h00000000;
		endcase
		
endmodule